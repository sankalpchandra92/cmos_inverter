magic
tech sky130A
timestamp 1753297477
<< nwell >>
rect -50 5 85 195
<< nmos >>
rect 10 -85 25 -40
<< pmos >>
rect 10 35 25 85
<< ndiff >>
rect -30 -50 10 -40
rect -30 -75 -20 -50
rect 0 -75 10 -50
rect -30 -85 10 -75
rect 25 -50 65 -40
rect 25 -75 35 -50
rect 55 -75 65 -50
rect 25 -85 65 -75
<< pdiff >>
rect -30 75 10 85
rect -30 50 -20 75
rect 0 50 10 75
rect -30 35 10 50
rect 25 70 65 85
rect 25 45 35 70
rect 55 45 65 70
rect 25 35 65 45
<< ndiffc >>
rect -20 -75 0 -50
rect 35 -75 55 -50
<< pdiffc >>
rect -20 50 0 75
rect 35 45 55 70
<< psubdiff >>
rect -30 -125 65 -115
rect -30 -145 -10 -125
rect 15 -145 65 -125
rect -30 -155 65 -145
<< nsubdiff >>
rect -30 160 65 170
rect -30 140 -10 160
rect 15 140 65 160
rect -30 130 65 140
<< psubdiffcont >>
rect -10 -145 15 -125
<< nsubdiffcont >>
rect -10 140 15 160
<< poly >>
rect 10 85 25 120
rect 10 20 25 35
rect -30 10 25 20
rect -30 -10 -20 10
rect 10 -10 25 10
rect -30 -20 25 -10
rect 10 -40 25 -20
rect 10 -100 25 -85
<< polycont >>
rect -20 -10 10 10
<< locali >>
rect -25 160 60 165
rect -25 140 -10 160
rect 15 140 60 160
rect -25 135 60 140
rect -25 85 5 135
rect -30 75 5 85
rect -30 50 -20 75
rect 0 50 5 75
rect -30 40 5 50
rect 30 70 65 80
rect 30 45 35 70
rect 55 45 65 70
rect 30 35 65 45
rect -30 10 10 20
rect -30 -10 -20 10
rect -30 -20 10 -10
rect 35 10 65 35
rect 35 -10 47 10
rect 35 -40 65 -10
rect -30 -50 5 -40
rect -30 -75 -20 -50
rect 0 -75 5 -50
rect -30 -85 5 -75
rect 30 -50 65 -40
rect 30 -75 35 -50
rect 55 -75 65 -50
rect 30 -85 65 -75
rect -25 -120 0 -85
rect -25 -125 60 -120
rect -25 -145 -10 -125
rect 15 -145 60 -125
rect -25 -150 60 -145
<< viali >>
rect -10 140 10 160
rect -20 -10 0 10
rect 47 -10 65 10
rect -10 -145 10 -125
<< metal1 >>
rect -105 160 20 165
rect -105 140 -10 160
rect 10 140 20 160
rect -105 135 20 140
rect -115 10 10 15
rect -115 -10 -20 10
rect 0 -10 10 10
rect -115 -15 10 -10
rect 40 10 165 15
rect 40 -10 47 10
rect 65 -10 165 10
rect 40 -15 165 -10
rect -100 -125 25 -120
rect -100 -145 -10 -125
rect 10 -145 25 -125
rect -100 -150 25 -145
<< labels >>
rlabel metal1 -95 145 -90 155 1 VDD
rlabel metal1 -92 -7 -87 3 1 VIN
rlabel metal1 114 -4 119 6 1 VOUT
rlabel metal1 -73 -141 -68 -131 1 GND
<< end >>
