** sch_path: /home/personal/Documents/inverter_folder/inverter1.sch
**.subckt inverter1
VDD VDD GND 1.8
VIN VIN GND 0
XM2 VOUT VIN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM1 VOUT VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
**** begin user architecture code
.lib /home/personal/pdk/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.dc VIN 0 1.8 0.01
.save all

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
